`timescale 1ns/1ns

module CA6_full_adder(input [7:0] A, B, output [7:0] result);
	assign result = A + B;	

endmodule