`timescale 1ns/1ns




module CA5_Q2_pre_synth(input clk, rst, j, output w);

	reg [2:0] ns, ps;
	parameter [2:0] A = 3'b000, B = 3'b001, C = 3'b010, D = 3'b011, E = 3'b100;

	always @(j, ps) begin

		ns <= 3'b0;
		
		case(ps)
		A: ns <= j ? B : A;
		B: ns <= j ? B : C;
		C: ns <= j ? B : D;
		D: ns <= j ? E : A;
		E: ns <= j ? B : C;
		default: ns <= 3'b0;
		endcase

	end

	assign w = (ps == E) ? ~j : 1'b0;



	always @(posedge clk, posedge rst) begin

		if (rst)
			ps <= 3'b0;
		else
			ps <= ns;





	end



endmodule